netcdf vgrid {
dimensions:
	nk = 50 ;
	nkp1 = 51 ;
variables:
	double dz(nk) ;
		dz:long_name = "z coordinate level thickness" ;
		dz:units = "m" ;
	double zt(nk) ;
		zt:long_name = "Diagnostic z coordinate level position" ;
		zt:comment = "Used for diagnostics only" ;
		zt:units = "m" ;
	double zw(nkp1) ;
		zw:long_name = "Diagnostic z coordinate interface position" ;
		zw:comment = "Used for diagnostics only" ;
		zw:units = "m" ;

// global attributes:
		:filename = "vgrid.nc" ;
data:

 dz = 10.1, 10.1, 10.1, 10.2, 10.2, 10.3, 10.5, 10.7, 10.9, 11.3, 11.7, 12.4, 
    13.3, 14.6, 16.3, 18.6, 21.7, 25.9, 31.4, 38.5, 47.4, 58.4, 71.3, 86, 
    101.9, 118.1, 134, 148.7, 161.6, 172.6, 181.5, 188.6, 194.1, 198.3, 
    201.4, 203.7, 205.4, 206.7, 207.6, 208.3, 208.7, 209.1, 209.3, 209.5, 
    209.7, 209.8, 209.8, 209.9, 209.9, 209 ;

 zt = 5.05, 15.15, 25.25, 35.4, 45.6, 55.85, 66.25, 76.85, 87.65, 98.75, 
    110.25, 122.3, 135.15, 149.1, 164.55, 182, 202.15, 225.95, 254.6, 289.55, 
    332.5, 385.4, 450.25, 528.9, 622.85, 732.85, 858.9, 1000.25, 1155.4, 
    1322.5, 1499.55, 1684.6, 1875.95, 2072.15, 2272, 2474.55, 2679.1, 
    2885.15, 3092.3, 3300.25, 3508.75, 3717.65, 3926.85, 4136.25, 4345.85, 
    4555.6, 4765.4, 4975.25, 5185.15, 5394.6 ;

 zw = 0, 10.1, 20.2, 30.3, 40.5, 50.7, 61, 71.5, 82.2, 93.1, 104.4, 116.1, 
    128.5, 141.8, 156.4, 172.7, 191.3, 213, 238.9, 270.3, 308.8, 356.2, 
    414.6, 485.9, 571.9, 673.8, 791.9, 925.9, 1074.6, 1236.2, 1408.8, 1590.3, 
    1778.9, 1973, 2171.3, 2372.7, 2576.4, 2781.8, 2988.5, 3196.1, 3404.4, 
    3613.1, 3822.2, 4031.5, 4241, 4450.7, 4660.5, 4870.3, 5080.2, 5290.1, 
    5499.1 ;
}
