netcdf vgrid {
dimensions:
	nz = 75 ;
	zt = 50 ;
	zw = 51 ;
variables:
	double dz(nz) ;
		dz:long_name = "z coordinate level thickness" ;
		dz:units = "m" ;
	double zt(zt) ;
		zt:long_name = "Diagnostic z coordinate level position" ;
		zt:comment = "Used for diagnostics only" ;
		zt:units = "m" ;
	double zw(zw) ;
		zw:long_name = "Diagnostic z coordinate interface position" ;
		zw:comment = "Used for diagnostics only" ;
		zw:units = "m" ;

// global attributes:
		:filename = "vgrid_cm4_10.nc" ;
data:

 dz = 10.00, 10.00, 10.00, 10.01, 10.02, 10.03, 10.05, 10.09, 10.13, 10.20, 10.29, 10.39, 10.53, 10.71, 10.91, 11.15, 11.46, 11.80, 12.22, 12.69, 13.24, 13.88, 14.62, 15.45, 16.40, 17.50, 18.72, 20.13, 21.70, 23.48, 25.47, 27.71, 30.22, 33.00, 36.08, 39.51, 43.26, 47.38, 51.86, 56.72, 61.95, 67.53, 73.47, 79.72, 86.25, 93.00, 99.95, 106.99, 114.09, 121.13, 128.08, 134.83, 141.32, 147.47, 153.23, 158.55, 163.40, 167.73, 171.57, 174.87, 177.70, 180.06, 181.97, 183.49, 184.66, 185.55, 186.17, 186.60, 186.87, 187.04, 187.11, 187.15, 187.16, 187.16, 187.17;

 zt = 5.05, 15.15, 25.25, 35.4, 45.6, 55.85, 66.25, 76.85, 87.65, 98.75, 
    110.25, 122.3, 135.15, 149.1, 164.55, 182, 202.15, 225.95, 254.6, 289.55, 
    332.5, 385.4, 450.25, 528.9, 622.85, 732.85, 858.9, 1000.25, 1155.4, 
    1322.5, 1499.55, 1684.6, 1875.95, 2072.15, 2272, 2474.55, 2679.1, 
    2885.15, 3092.3, 3300.25, 3508.75, 3717.65, 3926.85, 4136.25, 4345.85, 
    4555.6, 4765.4, 4975.25, 5185.15, 5394.6 ;

 zw = 0, 10.1, 20.2, 30.3, 40.5, 50.7, 61, 71.5, 82.2, 93.1, 104.4, 116.1, 
    128.5, 141.8, 156.4, 172.7, 191.3, 213, 238.9, 270.3, 308.8, 356.2, 
    414.6, 485.9, 571.9, 673.8, 791.9, 925.9, 1074.6, 1236.2, 1408.8, 1590.3, 
    1778.9, 1973, 2171.3, 2372.7, 2576.4, 2781.8, 2988.5, 3196.1, 3404.4, 
    3613.1, 3822.2, 4031.5, 4241, 4450.7, 4660.5, 4870.3, 5080.2, 5290.1, 
    5499.1 ;
}
