netcdf vgrid_75_2m {
dimensions:
	nz = 75 ;
	zt = 50 ;
	zw = 51 ;
variables:
	double dz(nz) ;
		dz:long_name = "z coordinate level thickness" ;
		dz:units = "m" ;
	double zt(zt) ;
		zt:long_name = "Diagnostic z coordinate level position" ;
		zt:comment = "Used for diagnostics only" ;
		zt:units = "m" ;
	double zw(zw) ;
		zw:long_name = "Diagnostic z coordinate interface position" ;
		zw:comment = "Used for diagnostics only" ;
		zw:units = "m" ;

// global attributes:
		:filename = "vgrid_75_2m.nc" ;
data:

 dz = 2, 2, 2, 2, 2.01, 2.01, 2.02, 2.03, 2.05, 2.08, 2.11, 2.15, 2.2, 2.27, 
    2.34, 2.44, 2.55, 2.69, 2.85, 3.04, 3.27, 3.54, 3.85, 4.22, 4.66, 5.18, 
    5.79, 6.52, 7.37, 8.37, 9.55, 10.94, 12.57, 14.48, 16.72, 19.33, 22.36, 
    25.87, 29.91, 34.53, 39.79, 45.72, 52.37, 59.76, 67.89, 76.74, 86.29, 
    96.47, 107.2, 118.35, 129.81, 141.42, 153.01, 164.41, 175.47, 186.01, 
    195.9, 205.01, 213.27, 220.6, 226.99, 232.43, 236.96, 240.63, 243.52, 
    245.72, 247.33, 248.45, 249.18, 249.62, 249.86, 249.96, 249.99, 250, 250 ;

 zt = 5.05, 15.15, 25.25, 35.4, 45.6, 55.85, 66.25, 76.85, 87.65, 98.75, 
    110.25, 122.3, 135.15, 149.1, 164.55, 182, 202.15, 225.95, 254.6, 289.55, 
    332.5, 385.4, 450.25, 528.9, 622.85, 732.85, 858.9, 1000.25, 1155.4, 
    1322.5, 1499.55, 1684.6, 1875.95, 2072.15, 2272, 2474.55, 2679.1, 
    2885.15, 3092.3, 3300.25, 3508.75, 3717.65, 3926.85, 4136.25, 4345.85, 
    4555.6, 4765.4, 4975.25, 5185.15, 5394.6 ;

 zw = 0, 10.1, 20.2, 30.3, 40.5, 50.7, 61, 71.5, 82.2, 93.1, 104.4, 116.1, 
    128.5, 141.8, 156.4, 172.7, 191.3, 213, 238.9, 270.3, 308.8, 356.2, 
    414.6, 485.9, 571.9, 673.8, 791.9, 925.9, 1074.6, 1236.2, 1408.8, 1590.3, 
    1778.9, 1973, 2171.3, 2372.7, 2576.4, 2781.8, 2988.5, 3196.1, 3404.4, 
    3613.1, 3822.2, 4031.5, 4241, 4450.7, 4660.5, 4870.3, 5080.2, 5290.1, 
    5499.1 ;
}
