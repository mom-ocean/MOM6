netcdf layer_coord {
dimensions:
	Layer = 75 ;
variables:
	double Layer(Layer) ;
		Layer:long_name = "Layer Target Potential Density" ;
		Layer:units = "kg m-3" ;

data:

 Layer =
    1009.420, 1012.893, 1016.366, 1019.839, 1023.311, 1026.784, 1030.169,
    1030.916, 1031.516, 1031.995, 1032.382, 1032.708, 1032.995, 1033.254,
    1033.497, 1033.729, 1033.950, 1034.162, 1034.366, 1034.558, 1034.740,
    1034.913, 1035.075, 1035.227, 1035.369, 1035.499, 1035.618, 1035.728,
    1035.829, 1035.922, 1036.009, 1036.089, 1036.164, 1036.234, 1036.301,
    1036.365, 1036.427, 1036.487, 1036.546, 1036.603, 1036.660, 1036.715,
    1036.768, 1036.815, 1036.856, 1036.893, 1036.926, 1036.955, 1036.981,
    1037.004, 1037.024, 1037.042, 1037.059, 1037.074, 1037.088, 1037.101,
    1037.115, 1037.128, 1037.142, 1037.155, 1037.168, 1037.182, 1037.195,
    1037.210, 1037.226, 1037.245, 1037.268, 1037.297, 1037.339, 1037.397,
    1037.468, 1037.558, 1037.665, 1037.783, 1037.900 ;
}
