netcdf layer_coord {
dimensions:
        Layer = 50 ;
variables:
        double Layer(Layer) ;

data:

 Layer = 1009.42, 1013.565, 1017.71, 1021.855, 1026, 1030.145, 1031.037,
    1031.719, 1032.229, 1032.633, 1032.978, 1033.288, 1033.575, 1033.846,
    1034.103, 1034.347, 1034.577, 1034.793, 1034.995, 1035.181, 1035.352,
    1035.507, 1035.648, 1035.776, 1035.891, 1035.996, 1036.092, 1036.181,
    1036.263, 1036.341, 1036.415, 1036.487, 1036.557, 1036.625, 1036.693,
    1036.757, 1036.814, 1036.863, 1036.905, 1036.943, 1036.975, 1037.003,
    1037.027, 1037.048, 1037.067, 1037.084, 1037.1, 1037.116, 1037.132,
    1037.148;
}
