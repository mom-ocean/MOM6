netcdf vgrid {
dimensions:
	nz = 75 ;
	zt = 50 ;
	zw = 51 ;
variables:
	double dz(nz) ;
		dz:long_name = "z coordinate level thickness" ;
		dz:units = "m" ;
	double zt(zt) ;
		zt:long_name = "Diagnostic z coordinate level position" ;
		zt:comment = "Used for diagnostics only" ;
		zt:units = "m" ;
	double zw(zw) ;
		zw:long_name = "Diagnostic z coordinate interface position" ;
		zw:comment = "Used for diagnostics only" ;
		zw:units = "m" ;

// global attributes:
		:filename = "vgrid_cm4_4.nc" ;
data:

 dz = 4.00, 4.00, 4.00, 4.00, 4.01, 4.02, 4.03, 4.05, 4.07, 4.11, 4.16, 4.22, 4.29, 4.39, 4.51, 4.65, 4.81, 5.02, 5.26, 5.54, 5.87, 6.26, 6.71, 7.24, 7.85, 8.57, 9.40, 10.36, 11.47, 12.76, 14.26, 15.97, 17.95, 20.22, 22.81, 25.79, 29.15, 32.95, 37.24, 42.02, 47.33, 53.20, 59.62, 66.57, 74.05, 82.03, 90.42, 99.17, 108.19, 117.37, 126.60, 135.76, 144.72, 153.37, 161.60, 169.30, 176.40, 182.82, 188.55, 193.56, 197.83, 201.44, 204.37, 206.72, 208.54, 209.90, 210.88, 211.54, 211.96, 212.22, 212.34, 212.40, 212.41, 212.41, 212.42;

 zt = 5.05, 15.15, 25.25, 35.4, 45.6, 55.85, 66.25, 76.85, 87.65, 98.75, 
    110.25, 122.3, 135.15, 149.1, 164.55, 182, 202.15, 225.95, 254.6, 289.55, 
    332.5, 385.4, 450.25, 528.9, 622.85, 732.85, 858.9, 1000.25, 1155.4, 
    1322.5, 1499.55, 1684.6, 1875.95, 2072.15, 2272, 2474.55, 2679.1, 
    2885.15, 3092.3, 3300.25, 3508.75, 3717.65, 3926.85, 4136.25, 4345.85, 
    4555.6, 4765.4, 4975.25, 5185.15, 5394.6 ;

 zw = 0, 10.1, 20.2, 30.3, 40.5, 50.7, 61, 71.5, 82.2, 93.1, 104.4, 116.1, 
    128.5, 141.8, 156.4, 172.7, 191.3, 213, 238.9, 270.3, 308.8, 356.2, 
    414.6, 485.9, 571.9, 673.8, 791.9, 925.9, 1074.6, 1236.2, 1408.8, 1590.3, 
    1778.9, 1973, 2171.3, 2372.7, 2576.4, 2781.8, 2988.5, 3196.1, 3404.4, 
    3613.1, 3822.2, 4031.5, 4241, 4450.7, 4660.5, 4870.3, 5080.2, 5290.1, 
    5499.1 ;
}
