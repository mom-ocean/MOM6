netcdf vgrid {
dimensions:
	nz = 75 ;
	zt = 50 ;
	zw = 51 ;
variables:
	double dz(nz) ;
		dz:long_name = "z coordinate level thickness" ;
		dz:units = "m" ;
	double zt(zt) ;
		zt:long_name = "Diagnostic z coordinate level position" ;
		zt:comment = "Used for diagnostics only" ;
		zt:units = "m" ;
	double zw(zw) ;
		zw:long_name = "Diagnostic z coordinate interface position" ;
		zw:comment = "Used for diagnostics only" ;
		zw:units = "m" ;

// global attributes:
		:filename = "vgrid_cm4.nc" ;
data:

 dz = 2.00, 2.00, 2.00, 2.00, 2.01, 2.01, 2.02, 2.02, 2.05, 2.07, 2.09, 2.13, 2.18, 2.24, 2.30, 2.40, 2.50, 2.62, 2.78, 2.95, 3.17, 3.42, 3.71, 4.07, 4.48, 4.97, 5.55, 6.23, 7.04, 7.99, 9.11, 10.43, 11.98, 13.80, 15.94, 18.42, 21.32, 24.66, 28.51, 32.91, 37.92, 43.56, 49.87, 56.88, 64.55, 72.91, 81.87, 91.40, 101.39, 111.73, 122.29, 132.93, 143.47, 153.78, 163.70, 173.07, 181.78, 189.76, 196.89, 203.17, 208.58, 213.14, 216.87, 219.87, 222.19, 223.94, 225.18, 226.04, 226.59, 226.90, 227.07, 227.14, 227.16, 227.16, 227.17;

 zt = 5.05, 15.15, 25.25, 35.4, 45.6, 55.85, 66.25, 76.85, 87.65, 98.75, 
    110.25, 122.3, 135.15, 149.1, 164.55, 182, 202.15, 225.95, 254.6, 289.55, 
    332.5, 385.4, 450.25, 528.9, 622.85, 732.85, 858.9, 1000.25, 1155.4, 
    1322.5, 1499.55, 1684.6, 1875.95, 2072.15, 2272, 2474.55, 2679.1, 
    2885.15, 3092.3, 3300.25, 3508.75, 3717.65, 3926.85, 4136.25, 4345.85, 
    4555.6, 4765.4, 4975.25, 5185.15, 5394.6 ;

 zw = 0, 10.1, 20.2, 30.3, 40.5, 50.7, 61, 71.5, 82.2, 93.1, 104.4, 116.1, 
    128.5, 141.8, 156.4, 172.7, 191.3, 213, 238.9, 270.3, 308.8, 356.2, 
    414.6, 485.9, 571.9, 673.8, 791.9, 925.9, 1074.6, 1236.2, 1408.8, 1590.3, 
    1778.9, 1973, 2171.3, 2372.7, 2576.4, 2781.8, 2988.5, 3196.1, 3404.4, 
    3613.1, 3822.2, 4031.5, 4241, 4450.7, 4660.5, 4870.3, 5080.2, 5290.1, 
    5499.1 ;
}
